module not_32bit(data_in, data_out);
    input [31:0] data_in;
    output [31:0] data_out;

    not NOT0(data_out[0], data_in[0]);
    not NOT1(data_out[1], data_in[1]);
    not NOT2(data_out[2], data_in[2]);
    not NOT3(data_out[3], data_in[3]);
    not NOT4(data_out[4], data_in[4]);
    not NOT5(data_out[5], data_in[5]);
    not NOT6(data_out[6], data_in[6]);
    not NOT7(data_out[7], data_in[7]);
    not NOT8(data_out[8], data_in[8]);
    not NOT9(data_out[9], data_in[9]);
    not NOT10(data_out[10], data_in[10]);
    not NOT11(data_out[11], data_in[11]);
    not NOT12(data_out[12], data_in[12]);
    not NOT13(data_out[13], data_in[13]);
    not NOT14(data_out[14], data_in[14]);
    not NOT15(data_out[15], data_in[15]);
    not NOT16(data_out[16], data_in[16]);
    not NOT17(data_out[17], data_in[17]);
    not NOT18(data_out[18], data_in[18]);
    not NOT19(data_out[19], data_in[19]);
    not NOT20(data_out[20], data_in[20]);
    not NOT21(data_out[21], data_in[21]);
    not NOT22(data_out[22], data_in[22]);
    not NOT23(data_out[23], data_in[23]);
    not NOT24(data_out[24], data_in[24]);
    not NOT25(data_out[25], data_in[25]);
    not NOT26(data_out[26], data_in[26]);
    not NOT27(data_out[27], data_in[27]);
    not NOT28(data_out[28], data_in[28]);
    not NOT29(data_out[29], data_in[29]);
    not NOT30(data_out[30], data_in[30]);
    not NOT31(data_out[31], data_in[31]);

endmodule